// module for calculating concentration
// modulate for calculating currents
