// may be more efficient to use fpga with arm processor on board
// to handle builtin ethernet traffic and move data to fpga
