// up to n preset spikes at preset positions then loop
