// specify inputs to a given node
// each node that can connect to another node has a signal
// if on, then that node is considered inputted
// could feed these inputs into an aggregator of sorts

// or could look at a crossbar impl

module matrix_flow(

);
endmodule
