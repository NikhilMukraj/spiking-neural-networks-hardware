// determine max number of numbers to store
// determine which operations to use (can be hardcoded and generated with eq hls)
// route correct numbers into operation
// store new numbers, potentially replacing old ones
// determine next operation
